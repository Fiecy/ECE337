// $Id: $
// File name:   sr_9bit.sv
// Created:     9/19/2016
// Author:      Yi Li
// Lab Section: 337-03
// Version:     1.0  Initial Design Entry
// Description: .
module sr_9bit
  (
   input 	clk,
   input 	n_rst,
   input 	shift_strobe,
   input 	serial_in,
   output [7:0] packet_data,
   output 	stop_bit
   );

   reg [8:0] 	p_out;

   flex_stp_sr #(.NUM_BITS(9), .SHIFT_MSB(0)) SHIFT(.clk(clk), .n_rst(n_rst), .shift_enable(shift_strobe), .serial_in(serial_in), .parallel_out(p_out));

   assign packet_data = p_out[7:0];
   assign stop_bit = p_out[8];

endmodule // sr_9bit
